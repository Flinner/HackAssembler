module main

type Symbols = map[string]int

fn init_symbols() Symbols {
	symbols := map{
		'__last_allocated__':  15// for allocating extra symbols
		'R0':  0
		'R1':  1
		'R2':  2
		'R3':  3
		'R4':  4
		'R5':  5
		'R6':  6
		'R7':  7
		'R8':  8
		'R9':  9
		'R10': 10
		'R11': 11
		'R12': 12
		'R13': 13
		'R14': 14
		'R15': 15
		'SP': 0
		'LCL': 1
		'ARG': 2
		'THIS': 3
		'THAT': 4
		'SCREEN': 16384
		'KBD': 24576
	}
	return symbols
}

fn (mut symbols Symbols) new(label string) int {
	a := symbols['__last_allocated__'] +1
	symbols[label]= a
	
	symbols['__last_allocated__'] = a
	return a
}

fn (mut symbols Symbols) write(label string, i int) {
	symbols[label] = i
}
