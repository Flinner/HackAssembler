module main

fn test_aa() {
	assert true
}

fn test_ab() {
	assert false
}
