module main

// tf! no way to convert ints to binary :|
// decbin converts to binary
fn decbin(n int) string {
	mut s := []string{len: 16, init: '0'}
	mut u := n

	for i := 0; u > 0; i++ {
		s[i] = if u & 1 == 1 { '1' } else { '0' }
		u = u >> 1
	}
	return s.join('').reverse()
}

// includes a field
const comp_map = map{
	'0':   '0101010'
	'1':   '0111111'
	'-1':  '0111010'
	'D':   '0001100'
	'A':   '0110000'
	'!D':  '0001101'
	'!A':  '0110001'
	'-D':  '0001111'
	'-A':  '0110011'
	'D+1': '0011111'
	'A+1': '0110111'
	'D-1': '0001110'
	'A-1': '0110010'
	'D+A': '0000010'
	'D-A': '0010011'
	'A-D': '0000111'
	'D&A': '0000000'
	'D|A': '0010101'
	'M':   '1110000'
	'!M':  '1110001'
	'-M':  '1110011'
	'M+1': '1110111'
	'M-1': '1110010'
	'D+M': '1000010'
	'D-M': '1010011'
	'M-D': '1000111'
	'D&M': '1000000'
	'D|M': '1010101'
}

const dest_map = map{
	'null': '000'
	'M':    '001'
	'D':    '010'
	'MD':   '011'
	'A':    '100'
	'AM':   '101'
	'AD':   '110'
	'AMD':  '111'
}

const jump_map = map{
	'null': '000'
	'JGT':  '001'
	'JEQ':  '010'
	'JGE':  '011'
	'JLT':  '100'
	'JNE':  '101'
	'JLE':  '110'
	'JMP':  '111'
}
