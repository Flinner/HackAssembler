module main

type Symbols = map[string]int

fn init_symbols() Symbols {
	symbols := map{
		'R0':  0
		'R1':  1
		'R2':  2
		'R3':  3
		'R4':  4
		'R5':  5
		'R6':  6
		'R7':  7
		'R8':  8
		'R9':  9
		'R10': 10
		'R11': 11
		'R12': 12
		'R13': 13
		'R14': 14
		'R15': 15
	}
	return symbols
}

fn (map Symbols) new(label string) int {
	return 99
}
