module main

fn main() {
	settings := handle_args()
}
